package agent_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "seq_item.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "sequencer.sv"
    `include "agent.sv"

    `include "sequence.sv"

endpackage
